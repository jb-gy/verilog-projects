module ORgate (a,b,y);

    input a,b;
    output y;