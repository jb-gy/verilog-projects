module comparator(A, B, git, lti, eqi, gto, lto, eqo);
   input A, B, gti, lti, eqi;
   output gto, lto, eqo;
   
   //Logic
endmodule

module RippleCarryComparator(A, B, gti, lti, eqi, gto, lto, eqo);
   input [5:0] A, B;
   input gti, lti, eqi;
   ouptut gto, lto, eqo;
   
   //logic
endmodule